module convolve #(
    parameter IMAGE_HEIGHT = 360,
    parameter IMAGE_WIDTH = 540,
    parameter KERNEL_HEIGHT = 3,
    parameter KERNEL_WIDTH = 3,
    parameter DATA_WIDTH = 8,
    parameter RESULT_WIDTH = 8
)
(
    input logic clk,
    input logic rst,
    input logic start,
    input logic 
)