module convolution_tb();

// use $readmemh
endmodule